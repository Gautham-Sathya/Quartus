LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

entity 4bCounter is port (                 	
   CP: 	in std_logic; 	-- clock
   SR:  in std_logic;  -- Active low, synchronous reset
   P:    in std_logic_vector(3 downto 0);  -- Parallel input
   PE:   in std_logic;  -- Parallel Enable (Load)
   CEP: in std_logic;  -- Count enable parallel input
   CET:  in std_logic; -- Count enable trickle input
   Q:   out std_logic_vector(3 downto 0);            			
    TC:  out std_logic  -- Terminal Count
);            		
end 4bCounter;

architecture model of 4bCounter is
signal Q_in: std_logic_vector(3 downto 0);
begin

process ( CP)
begin
if(rising_edge(CP)) then
	if SR = '0' then  Q_in <= "0000";
	elsif PE = '1' then Q_in<=P;
	elsif CEP = '1' and CET = '1' then Q_in<= std_logic_vector(unsigned(Q_in)+1);
	end if;

end if;


end process;
Q <= Q_in;
TC<= Q_in(0) and Q_in(1) and Q_in(2) and Q_in(3);

end model;
